module Full_Adder_3_bit (
    input  logic [2:0] A,
    input  logic [2:0] B,
    output logic [3:0] Sum
);
    logic c1, c2;

    Full_Adder FA0 (.A(A[0]), .B(B[0]), .Cin(1'b0), .Sum(Sum[0]), .Cout(c1));
    Full_Adder FA1 (.A(A[1]), .B(B[1]), .Cin(c1),   .Sum(Sum[1]), .Cout(c2));
    Full_Adder FA2 (.A(A[2]), .B(B[2]), .Cin(c2),   .Sum(Sum[2]), .Cout(Sum[3]));
endmodule
